module spem
    (
    input wire [3:0] data_in,
    output wire [3:0] data_out
    );



endmodule: spem