module aes_core
    (
    input logic clk,
	input logic rst,
    input logic [127:0] data_in,
    input logic [127:0] round_key,
    output logic [127:0] data_out
    );



endmodule: aes_core
